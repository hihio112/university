`timescale 1ns / 1ps

module tb_dct();
reg clk;
reg rst_n;
reg signed [7:0] x[0:7][0:7];
wire signed [19:0] Y[0:7][0:7];
wire r_vaild;

integer i = 0;
integer j = 0;
integer fd;
always #5 clk = ~clk;   // T = 10ns

initial begin
    fd = $fopen("my_file.txt", "w");  
    clk = 0;
    rst_n = 0;
    $srandom(1);
    
    for(i=0;i<8;i=i+1) begin
        for(j=0;j<8;j=j+1) begin
            x[i][j] = $random%256;
            $fwrite(fd, x[i][j]); 
            end
         $fwrite(fd, "\n"); 
         end
    #10 rst_n = 1;
    $fclose(fd);
    #2000 $finish;
end

dct_1d_full
#(
   .N(8)
) tb_full_dct
(
.clk(clk),
.rst_n(rst_n),
//zero row
.x00(x[0][0]), 
.x01(x[0][1]),
.x02(x[0][2]),
.x03(x[0][3]),
.x04(x[0][4]),
.x05(x[0][5]),
.x06(x[0][6]),
.x07(x[0][7]),
.x10(x[1][0]),
.x11(x[1][1]),
.x12(x[1][2]),
.x13(x[1][3]),
.x14(x[1][4]),
.x15(x[1][5]),
.x16(x[1][6]),
.x17(x[1][7]),
.x20(x[2][0]),
.x21(x[2][1]),
.x22(x[2][2]),
.x23(x[2][3]),
.x24(x[2][4]),
.x25(x[2][5]),
.x26(x[2][6]),
.x27(x[2][7]),
.x30(x[3][0]),
.x31(x[3][1]),
.x32(x[3][2]),
.x33(x[3][3]),
.x34(x[3][4]),
.x35(x[3][5]),
.x36(x[3][6]),
.x37(x[3][7]),
.x40(x[4][0]),
.x41(x[4][1]),
.x42(x[4][2]),
.x43(x[4][3]),
.x44(x[4][4]),
.x45(x[4][5]),
.x46(x[4][6]),
.x47(x[4][7]),
.x50(x[5][0]),
.x51(x[5][1]),
.x52(x[5][2]),
.x53(x[5][3]),
.x54(x[5][4]),
.x55(x[5][5]),
.x56(x[5][6]),
.x57(x[5][7]),
.x60(x[4][0]),
.x61(x[6][1]),
.x62(x[6][2]),
.x63(x[6][3]),
.x64(x[6][4]),
.x65(x[6][5]),
.x66(x[6][6]),
.x67(x[6][7]),
.x70(x[7][0]),
.x71(x[7][1]),
.x72(x[7][2]),
.x73(x[7][3]),
.x74(x[7][4]),
.x75(x[7][5]),
.x76(x[7][6]),
.x77(x[7][7]),
.Y00(Y[0][0]), 
.Y01(Y[0][1]),
.Y02(Y[0][2]),
.Y03(Y[0][3]),
.Y04(Y[0][4]),
.Y05(Y[0][5]),
.Y06(Y[0][6]),
.Y07(Y[0][7]),
.Y10(Y[1][0]),
.Y11(Y[1][1]),
.Y12(Y[1][2]),
.Y13(Y[1][3]),
.Y14(Y[1][4]),
.Y15(Y[1][5]),
.Y16(Y[1][6]),
.Y17(Y[1][7]),
.Y20(Y[2][0]),
.Y21(Y[2][1]),
.Y22(Y[2][2]),
.Y23(Y[2][3]),
.Y24(Y[2][4]),
.Y25(Y[2][5]),
.Y26(Y[2][6]),
.Y27(Y[2][7]),
.Y30(Y[3][0]),
.Y31(Y[3][1]),
.Y32(Y[3][2]),
.Y33(Y[3][3]),
.Y34(Y[3][4]),
.Y35(Y[3][5]),
.Y36(Y[3][6]),
.Y37(Y[3][7]),
.Y40(Y[4][0]),
.Y41(Y[4][1]),
.Y42(Y[4][2]),
.Y43(Y[4][3]),
.Y44(Y[4][4]),
.Y45(Y[4][5]),
.Y46(Y[4][6]),
.Y47(Y[4][7]),
.Y50(Y[5][0]),
.Y51(Y[5][1]),
.Y52(Y[5][2]),
.Y53(Y[5][3]),
.Y54(Y[5][4]),
.Y55(Y[5][5]),
.Y56(Y[5][6]),
.Y57(Y[5][7]),
.Y60(Y[6][0]),
.Y61(Y[6][1]),
.Y62(Y[6][2]),
.Y63(Y[6][3]),
.Y64(Y[6][4]),
.Y65(Y[6][5]),
.Y66(Y[6][6]),
.Y67(Y[6][7]),
.Y70(Y[7][0]),
.Y71(Y[7][1]),
.Y72(Y[7][2]),
.Y73(Y[7][3]),
.Y74(Y[7][4]),
.Y75(Y[7][5]),
.Y76(Y[7][6]),
.Y77(Y[7][7])
);
endmodule
